/** @copyright (C) 2018,  Gavin J Stark.  All rights reserved.
 *
 * @copyright
 *    Licensed under the Apache License, Version 2.0 (the "License");
 *    you may not use this file except in compliance with the License.
 *    You may obtain a copy of the License at
 *     http://www.apache.org/licenses/LICENSE-2.0.
 *   Unless required by applicable law or agreed to in writing, software
 *   distributed under the License is distributed on an "AS IS" BASIS,
 *   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 *   See the License for the specific language governing permissions and
 *   limitations under the License.
 *
 * @file   tb_riscv_minimal.cdl
 * @brief  Testbench for minimal RISC-V
 *
 */

/*a Includes
 */
include "apb::apb.h"
include "apb::apb_targets.h"
include "jtag.h"
include "jtag_modules.h"

/*a External modules
extern module se_test_harness( clock clk, output t_jtag jtag, output bit tck_enable, input bit tdo )
{
    timing from rising clock clk jtag, tck_enable;
    timing to rising clock clk tdo;
}
 */
/*a Module
 */
module tb_jtag_apb_timer( clock jtag_tck, // Test harness runs off this
                          clock apb_clock,
                          input bit reset_n,
                          input  t_apb_request  apb_request  "APB request",
                          output t_apb_response apb_response "APB response",
                          input bit tck_enable "Clock enable for actual JTAG clock",
                          input t_jtag jtag,
                          output bit tdo
)
{

    /*b Nets
     */
    net t_apb_response apb_response;
    net t_jtag apb_jtag;
    net bit apb_jtag_tck_enable;
    comb t_jtag jtag_int;
    net bit tdo;
    net bit[5]ir;
    net t_jtag_action dr_action;
    net bit[50]dr_in;
    net bit[50]dr_tdi_mask;
    net bit[50]dr_out;
    net t_apb_request apb_request_int;
    net t_apb_response apb_response_int;
    net bit[3] timer_equalled;
    comb bit tck_enable_fix;
    gated_clock clock jtag_tck active_high tck_enable_fix jtag_tck_gated;

    /*b Instantiate APB timer
     */
    dut_instance: {
        tck_enable_fix = tck_enable | apb_jtag_tck_enable;
        apb_target_jtag apb2jtag( clk <- jtag_tck,
                                  reset_n <= reset_n,

                                  apb_request <= apb_request,
                                  apb_response => apb_response,
                                  jtag_tck_enable => apb_jtag_tck_enable,
                                  jtag => apb_jtag,
                                  jtag_tdo <= tdo
            );
        jtag_int  = jtag;
        jtag_int |= apb_jtag;
        jtag_tap tap( jtag_tck <- jtag_tck_gated,
                      reset_n <= reset_n,
                      jtag <= jtag_int,
                      tdo => tdo,

                      ir => ir,
                      dr_action => dr_action,
                      dr_in => dr_in,
                      dr_tdi_mask <= dr_tdi_mask,
                      dr_out <= dr_out );

        jtag_tap_apb apb( jtag_tck <- jtag_tck_gated,
                      reset_n <= reset_n,

                      ir <= ir,
                      dr_action <= dr_action,
                      dr_in <= dr_in,
                      dr_tdi_mask => dr_tdi_mask,
                      dr_out => dr_out,

                      apb_clock <- apb_clock,
                      apb_request => apb_request_int,
                      apb_response <= apb_response_int );

        apb_target_timer timer( clk <- apb_clock,
                         reset_n <= reset_n,

                         apb_request <= apb_request_int,
                         apb_response => apb_response_int,

                         timer_equalled => timer_equalled
            );
    }
}
